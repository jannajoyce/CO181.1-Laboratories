`timescale 1ns / 1ps

/*
** -------------------------------------------------------------------
**  Instruction Rom for Single-Cycle MIPS Processor for Altera FPGAs
**
**  Change Log:
**  1/13/2012 - Adrian Caulfield - Initial Implementation
**
**
**  NOTE:  The Provided Modules do NOT follow the course coding standards
*/

module inst_rom (
	input	clock,
	input reset,
	input [31:0] addr_in, 
	output reg [31:0] data_out
);
	parameter ADDR_WIDTH = 5;
	//parameter INIT_PROGRAM="C:/intelFPGA_lite/18.1/quartus/181.1/lab6_jumao-as/quartus/blank.memh";
	parameter INIT_PROGRAM="C:/intelFPGA_lite/18.1/quartus/181.1/lab7_jumao-as/nbhelloworld.inst_rom.memh";

	reg [31:0] rom [0:(2**ADDR_WIDTH)-1];
	//reg [31:0] out;
	
	//assign data_out = {out[7:0],out[15:8],out[23:16],out[31:24]}; //flip bytes
	
	initial
	begin
		$readmemh(INIT_PROGRAM, rom);
	end
	
	always @(*) begin
		if (reset) begin
			data_out = 32'h00000000;
		end else begin
			data_out = {
                rom[addr_in[ADDR_WIDTH+1:2]][7:0], 
                rom[addr_in[ADDR_WIDTH+1:2]][15:8], 
                rom[addr_in[ADDR_WIDTH+1:2]][23:16], 
                rom[addr_in[ADDR_WIDTH+1:2]][31:24]
            };
        end
	end

endmodule

